// somewhat contrived, but i came across a real-life file that caused this
// crash.
value=
hello/
world;

// dummy stuff to generate a tag
module dummy;
endmodule
